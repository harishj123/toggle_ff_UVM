interface tff_interface(input logic clk);
  logic rstn;
  logic t;
  logic q;
endinterface
